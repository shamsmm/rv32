module cu(input logic [6:0] opcode);

endmodule