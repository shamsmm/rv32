// Connect to RV core

module clint (
    output bit irq_sw = 1'b0,
    output bit irq_ext = 1'b0,
    output bit irq_timer = 1'b0
);
    
endmodule